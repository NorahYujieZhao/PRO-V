
module RefModule (
  input a,
  input b,
  output q
);

  assign q = a&b;

endmodule
