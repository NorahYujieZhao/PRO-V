module top_module(
	input clk,
	input load,
	input [255:0] data,
	output reg [255:0] q);
	
	
	logic [323:0] q_pad;
	always@(*) begin
		for (int i=0;i<16;i++)
			q_pad[18*(i+1)+1 +: 16] = q[16*i +: 16];
		q_pad[1 +: 16] = q[16*15 +: 16];
		q_pad[18*17+1 +: 16] = q[0 +: 16];
		
		for (int i=0; i<18; i++) begin
			q_pad[i*18] = q_pad[i*18+16];
			q_pad[i*18+17] = q_pad[i*18+1];
		end
	end
	
	always @(posedge clk) begin
		for (int i=0;i<16;i++)
		for (int j=0;j<16;j++) begin
			q[i*16+j] <= 
				((q_pad[(i+1)*18+j+1 -1+18] + q_pad[(i+1)*18+j+1 +18] + q_pad[(i+1)*18+j+1 +1+18] +
				q_pad[(i+1)*18+j+1 -1]                                + q_pad[(i+1)*18+j+1+1] +
				q_pad[(i+1)*18+j+1 -1-18]   + q_pad[(i+1)*18+j+1 -18] + q_pad[(i+1)*18+j+1 +1-18]) & 3'h7 | q[i*16+j]) == 3'h3;
		end
		
		if (load)
			q <= data;
		
	end
	
endmodule
